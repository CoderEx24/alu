`include "alu.v"

module t_arthmetic_unit;
	reg [10: 0] in;
	wire [4: 0] result;
	wire C_out;

	arithmetic_unit
endmodule
